-- Averager

-- This module should take in an 8 bit input signal, a Sampling Clock Signal
-- (Goes high for 1 clock cycle (e.g. using a Safe Rising Edge component) when
-- a sample is taken from the ADC) and a master Clock Signal. It should read
-- the input signal on the rising edge of the clock when the Sampling Clock
-- Signal is high and then output the value of the input.

-- This module stores the last 4 input signals and adds them it then divides 
-- sum of the last 4 inputs by 4 and ouputs this - i.e. the average of the 
-- last 4 input signals

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


  
entity Averager is
  generic ( -- defines most of the constants defining filter behaviour
    -- Notation note: _1 = -1
    NoOfInputBits : integer := N1;
    NoOfInputBits_1 : integer := N2;
    DoubleNoOfInputBits_1 : integer := N3;
    NoOfBitsToShift : integer := N4;
    NoOfBitsToShift_1 : integer := N5;
    NoOfCoefs_1 : integer := N6;
    NoOfBitsForSumRegister : integer := N7;
    NoOfBitsForSumRegister_1 : integer := N8
  );

  port (
    clk : in std_logic;
    ClockEnable : in std_logic;
    Averager_In : in std_logic_vector(NoOfInputBits_1 downto 0);
    Averager_Out : out std_logic_vector(NoOfInputBits_1 downto 0)
    );
end Averager;

architecture AveragerArchitecture of Averager is
  type array_of_Nbit is array (0 to NoOfCoefs_1) of std_logic_vector(NoOfInputBits_1 downto 0);
  type array_of_2Nbit is array (0 to NoOfCoefs_1) of std_logic_vector(DoubleNoOfInputBits_1 downto 0);
  type array_N_integer is array (0 to NoOfCoefs_1) of integer;
  
  function "*"(a, b : array_of_Nbit) return array_of_2Nbit is
    variable result_v : array_of_2Nbit;
  begin
    for idx in result_v'range loop
      result_v(idx) := std_logic_vector(unsigned(a(idx)) * unsigned(b(idx)));
    end loop;
    return result_v;
  end function;

  function to_array_of_Nbit(v : array_N_integer; N : integer) return array_of_Nbit is
    variable result_v : array_of_Nbit;
  begin
    for idx in result_v'range loop
      result_v(idx) := std_logic_vector(to_unsigned(v(idx), N));
    end loop;
    return result_v;
  end function;

  -- signal and constant decleration
  constant Coefficients : array_of_Nbit := to_array_of_Nbit(N9, NoOfInputBits);
-- coefficients are defined on last line
  constant ZerosArray : std_logic_vector(NoOfBitsToShift_1 downto 0) := "N10";
  signal Array_Last4Vals : array_of_Nbit;
  --signal SumOfSignals : unsigned(7 downto 0); 
  signal ProductArray : array_of_2Nbit;
  signal SumOfSignals : std_logic_vector(NoOfBitsForSumRegister_1 downto 0);
  signal Average16Bits : std_logic_vector(NoOfBitsForSumRegister_1 downto 0);
begin
  process(clk, ClockEnable) is
  begin
--    report "working";
    if (rising_edge(clk) and ClockEnable = '1') then -- read in state when 
      -- ADC clock is high and master clock rises
--      report "read in :" & integer'image(to_integer(unsigned(Averager_In)));
      for i in NoOfCoefs_1 downto 1 loop
        Array_Last4Vals(i) <= Array_Last4Vals(i-1);
      end loop;
      Array_Last4Vals(0) <= Averager_In;
    end if;
    if (rising_edge(clk)) then
      ProductArray <= Coefficients*Array_Last4Vals;
      SumOfSignals <= std_logic_vector(to_unsigned(
        ADDITION_STUFF_GOES_HERE
        , NoOfBitsForSumRegister));
      Average16Bits <= ZerosArray & SumOfSignals(NoOfBitsForSumRegister_1 downto NoOfBitsToShift); -- divide by 2**NoOfBitsToShift (bitshift right by NoOfBitsToShift)
      Averager_Out <= Average16Bits(NoOfInputBits_1 downto 0); -- take 8 least significant bits
    end if;
  end process;
end AveragerArchitecture;
